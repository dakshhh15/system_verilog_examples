interface int1 (input logic clk, rst);
  logic d, q;
endinterface
