interface int1;
  logic a, b, sel, out;
endinterface
