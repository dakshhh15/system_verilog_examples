interface int1 (input logic clk, rst);
  logic [3:0] a, b;
  logic [4:0] sum;
  logic valid;
endinterface
