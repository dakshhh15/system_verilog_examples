interface int1;
  logic [3:0] sum, a, b;
  logic cin, cout;
endinterface
