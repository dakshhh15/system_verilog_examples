interface int1 (input logic clk, clr);
  logic [3:0] q, d;
  logic [1:0] s;
  logic sl, sr;
endinterface
