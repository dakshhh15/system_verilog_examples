//  https://verifasttechpvtltd-my.sharepoint.com/:x:/r/personal/vdoshi_verifasttech_com/_layouts/15/Doc.aspx?sourcedoc=%7B448A0860-E56C-4583-8532-3E4A71569FA5%7D&file=Internship%20_Tracker.xlsx&fromShare=true&action=default&mobileredirect=true
