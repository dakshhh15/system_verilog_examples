interface int1;
  logic [3:0] a, b, sum;
  logic cin, cout;
endinterface
