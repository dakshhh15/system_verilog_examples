interface int1 ();
  
  logic a, b, cin, carry, sum;
  
endinterface
